package tbArchPkg;
    import VtbPkg::*;
    import typesPkg::*;
    import scenarioPkg::*;
    import utilityPkg::*;
    import jobsPkg::*;
    `include "taskFactory.sv"
    `include "taskManager.sv"
    `include "scenarioGen.sv"
endpackage
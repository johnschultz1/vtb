package VtbPkg;
    import scenarioPkg::*;
    import typesPkg::*;
    import utilityPkg::*;
    `include "messageQ.sv"
endpackage
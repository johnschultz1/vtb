module dut(
    input clk,
    input rst
);
endmodule
package jobsPkg;

    `include "jobUtil.sv";
    `include "helloHuman.sv";

endpackage
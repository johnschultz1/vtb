package utilityPkg;
    import typesPkg::*;
    `include "utility.sv"
endpackage
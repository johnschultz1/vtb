package jobsPkg;
    import utilityPkg::*;

    `include "jobUtil.sv";
    `include "toggleSeq.sv";
    `include "helloHuman.sv";
    `include "inOrderScoreBoard.sv"
    `include "monitor.sv"
    `include "predictor.sv"
    `include "receiver.sv"
    `include "broadcaster.sv"
    `include "delay.sv"
    `include "dataGen.sv"
    `include "driver.sv"

endpackage
package jobsPkg;

    `include "jobUtil.sv";
    `include "toggleSeq.sv";
    `include "helloHuman.sv";

endpackage
package tbArchPkg;
    import VtbPkg::*;
    import typesPkg::*;
    import scenarioPkg::*;
    import utilityPkg::*;
    import jobsPkg::*;
    `include "jobFactory.sv"
    `include "jobManager.sv"
    `include "scenarioGen.sv"
endpackage
class delay;

    `startJob
        #(cfg.ints["CYCLES"]);
    `endJob

endclass;